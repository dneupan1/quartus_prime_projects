-- Lab4PartII 

-- Students
--		Deepak Neupane
--		Hansen Shamoon
--
-- In this lab, we are to implement an alternative way to specify a counter
-- by using a register and adding 1 to it's value. 
-- 		Q <= Q + 1  (incrementing register value as counter)

LIBRARY IEEE;
