--Lab Three Part III

--Students:
--	Hansen Shamoon 
--	Deepak Neupane

-- 
--

LIBRARY ieee;
USE ieee.std_logic_1164.all;


ENTITY LabThreePartIII is
    PORT ( 
				);
END LabThreePartIII;

ARCHITECTURE Behavior of LabThreePartII is


BEGIN 
	
END Behavior;
