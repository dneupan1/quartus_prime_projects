-- LabFourPartI
--
-- Students:
-- 	Deepak Neupane
--		Hansen Shamoon
--
-- In this part, we need to implement a 8 bit counter using 8 instances of 
-- T-Type flip flop

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.all;

