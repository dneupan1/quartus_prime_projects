-- Final Project
--
-- Students:
--	 Hansen Shamoon 
--	 Deepak Neupane
--  Digvijay Jonna
--
--


LIBRARY ieee;
USE ieee.std_logic_1164.all;

-- Four Bit Adder (Top Level Entity)
ENTITY FinalProject is
    PORT ( 
	 
	 );
END FinalProject;

ARCHITECTURE Behavioral of FinalProject is


BEGIN
	
    
END Behavioral;

